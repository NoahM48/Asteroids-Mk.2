module sevenSeg(a1, b1, c1, d1, a2, b2, c2, d2, a3, b3, c3, d3, a4, b4, c4, d4, o1, o2, o3, o4, o5, o6, o7, o12, o22, o32, o42, o52, o62, o72, o13, o23, o33, o43, o53, o63, o73, o14, o24, o34, o44, o54, o64, o74);

input a1, b1, c1, d1, a2, b2, c2, d2, a3, b3, c3, d3, a4, b4, c4, d4;
output o1, o2, o3, o4, o5, o6, o7, o12, o22, o32, o42, o52, o62, o72, o13, o23, o33, o43, o53, o63, o73, o14, o24, o34, o44, o54, o64, o74;

assign o1 = ~((~b1&&~d1) || (~a1&&c1) || (b1&&c1) || (a1&&~d1) || (~a1&&b1&&d1) || (a1&&~b1&&~c1));

assign o2 = ~((~a1&&~b1) || (~b1&&~d1) || (~a1&&~c1&&~d1) || (~a1&&c1&&d1) || (a1&&~c1&&d1));

assign o3 = ~((~a1&&~c1) || (~a1&&d1) || (~c1&&d1) || (~a1&&b1) || (a1&&~b1));

assign o4 = ~((~a1&&~b1&&~d1) || (~b1&&c1&&d1) || (b1&&~c1&&d1) || (b1&&c1&&~d1) || (a1&&~c1&&~d1));

assign o5 = ~((~b1&&~d1) || (c1&&~d1) || (a1&&c1) || (a1&&b1));

assign o6 = ~((~c1&&~d1) || (b1&&~d1) || (a1&&~b1) || (a1&&c1) || (~a1&&b1&&~c1));

assign o7 = ~((~b1&&c1) || (c1&&~d1) || (a1&&~b1) || (a1&&d1) || (~a1&&b1&&~c1));

assign o12 = ~((~b2&&~d2) || (~a2&&c2) || (b2&&c2) || (a2&&~d2) || (~a2&&b2&&d2) || (a2&&~b2&&~c2));

assign o22 = ~((~a2&&~b2) || (~b2&&~d2) || (~a2&&~c2&&~d2) || (~a2&&c2&&d2) || (a2&&~c2&&d2));

assign o32 = ~((~a2&&~c2) || (~a2&&d2) || (~c2&&d2) || (~a2&&b2) || (a2&&~b2));

assign o42 = ~((~a2&&~b2&&~d2) || (~b2&&c2&&d2) || (b2&&~c2&&d2) || (b2&&c2&&~d2) || (a2&&~c2&&~d2));

assign o52 = ~((~b2&&~d2) || (c2&&~d2) || (a2&&c2) || (a2&&b2));

assign o62 = ~((~c2&&~d2) || (b2&&~d2) || (a2&&~b2) || (a2&&c2) || (~a2&&b2&&~c2));

assign o72 = ~((~b2&&c2) || (c2&&~d2) || (a2&&~b2) || (a2&&d2) || (~a2&&b2&&~c2));

assign o13 = ~((~b3&&~d3) || (~a3&&c3) || (b3&&c3) || (a3&&~d3) || (~a3&&b3&&d3) || (a3&&~b3&&~c3));

assign o23 = ~((~a3&&~b3) || (~b3&&~d3) || (~a3&&~c3&&~d3) || (~a3&&c3&&d3) || (a3&&~c3&&d3));

assign o33 = ~((~a3&&~c3) || (~a3&&d3) || (~c3&&d3) || (~a3&&b3) || (a3&&~b3));

assign o43 = ~((~a3&&~b3&&~d3) || (~b3&&c3&&d3) || (b3&&~c3&&d3) || (b3&&c3&&~d3) || (a3&&~c3&&~d3));

assign o53 = ~((~b3&&~d3) || (c3&&~d3) || (a3&&c3) || (a3&&b3));

assign o63 = ~((~c3&&~d3) || (b3&&~d3) || (a3&&~b3) || (a3&&c3) || (~a3&&b3&&~c3));

assign o73 = ~((~b3&&c3) || (c3&&~d3) || (a3&&~b3) || (a3&&d3) || (~a3&&b3&&~c3));

assign o14 = ~((~b4&&~d4) || (~a4&&c4) || (b4&&c4) || (a4&&~d4) || (~a4&&b4&&d4) || (a4&&~b4&&~c4));

assign o24 = ~((~a4&&~b4) || (~b4&&~d4) || (~a4&&~c4&&~d4) || (~a4&&c4&&d4) || (a4&&~c4&&d4));

assign o34 = ~((~a4&&~c4) || (~a4&&d4) || (~c4&&d4) || (~a4&&b4) || (a4&&~b4));

assign o44 = ~((~a4&&~b4&&~d4) || (~b4&&c4&&d4) || (b4&&~c4&&d4) || (b4&&c4&&~d4) || (a4&&~c4&&~d4));

assign o54 = ~((~b4&&~d4) || (c4&&~d4) || (a4&&c4) || (a4&&b4));

assign o64 = ~((~c4&&~d4) || (b4&&~d4) || (a4&&~b4) || (a4&&c4) || (~a4&&b4&&~c4));

assign o74 =~((~b4&c4) | (c4&~d4) | (a4&~b4) | (a4&d4) | (~a4&b4&~c4));




endmodule